*** FACET 2X1-LAYOUT FROM LIBRARY GENNUMFLAT.ELIB ***
*** FACET CREATED MON OCT 08 14:34:20 2012
*** VERSION 1 LAST REVISED MON OCT 08 14:34:20 2012
*** EXTRACTED BY ELECTRIC DESIGN SYSTEM, VERSION 5.5.2
*** UC SPICE *** , MIN_RESIST 0.000000, MIN_CAPAC 0.000000FF
.OPTIONS NOMOD NOPAGE
*---------------------------------------------------------------------
* NOMINAL model set for GA911 semicustom array.  V1.1 July 1990
* Set 8 : NPR = NNN

.MODEL SNPN_911 NPN (IS=5E-17 BF=147 VAF=80 IKF=4.3E-3 ISE=8E-18 NE=1.233
+BR=1.9 VAR=11 IKR=6E-4 ISC=5E-16 NC=1.08 RE=12 RB=1200 RBM=200 RC=25
+CJE=58E-15 VJE=0.83 MJE=0.35 CJC=133E-15 VJC=0.6 MJC=0.44 XCJC=1
+CJS=830E-15 VJS=0.6 MJS=0.4 ISS=1E-16 FC=0.85 TF=60P XTF=48 ITF=3E-2
+TR=10N EG=1.16 XTI=3 XTB=1.6)

.MODEL LNPN_911 NPN (IS=7.5E-16 BF=206 VAF=58 IKF=20E-3 ISE=8E-18 NE=1.105
+BR=4.5 VAR=11 IKR=2E-3 NC=2 RE=0.7 RB=660 RBM=35 RC=9 CJE=550E-15 VJE=0.83
+MJE=0.35 CJC=440E-15 VJC=0.6 MJC=0.44 XCJC=1 CJS=1.65E-12 VJS= 0.6 MJS=0.4
+ISS=2E-16 FC=0.85 TF=70P XTF=20 ITF=0.2 TR=2N EG=1.16 XTI=3 XTB=1.6)

.MODEL CAP_NPN NPN (IS=10E-15 XTI=3 EG=1.16 VAF=31 BF=350 NE=1.45 ISE=1E-15
+IKF=0.5 XTB=1.6 BR=10 NC=2 RC=50 RB=1100 RBM=300 CJC=3.29E-12 MJC=0.44
+VJC=0.6 FC=0.85 CJE=8.8E-12 MJE=0.35 VJE=0.83 TR=10N TF=80E-12 ITF= 0.3 VTF=6
+XTF=50 CJS=3.27E-12 MJS=0.4 VJS=0.6 ISS=4E-16)

.MODEL JP90K PJF (VTO=-2.65 BETA=2.3E-6 BETATCE=-0.3 IS=1.8E-16 RS=650
+RD=3.5E3 CGD=250E-15 CGS=135E-15 M=0.38 PB=0.75)

.MODEL SPNP_911 LPNP (IS=2.9E-16 XTI=3.3 EG=1.16 VAF=60 BF=49 NE=1.585
+ISE=4E-15 IKF=140E-6 XTB=1.5 BR=0.5108 VAR=6 NC=1.58 ISC=40E-15 IKR=140E-6
+RC=50 RE=20 RB=150 RBM=30 CJC=245E-15 MJC=0.44 VJC=0.6 FC=0.85 CJE=54E-15
+MJE=0.44 VJE=0.6 TF=14E-9 ITF=3E-3 VTF=4 XTF=0.8 TR=338E-9
+ISS=1E-16 CJS=830E-15 VJS=0.6 MJS=0.4)

.MODEL SUB_PNP PNP (IS=8E-15 XTI=3.3 EG=1.16 VAF=100 BF=40 NE=1.49 ISE=35E-15
+IKF=4E-3 XTB=1.5 BR=.2 VAR=20 NC=2 RE=50 RC=70 RB=200 RBM=20 CJC=3.27E-12
+MJC=0.4 VJC=0.6 FC=0.85 CJE=3.29E-12 MJE=0.44 VJE=0.6 TR=633E-9 TF=10E-9
+ITF=30E-3 VTF=50 XTF=1.2)

.MODEL RP- RES (R=1.0 TC1=1.12E-3 TC2=2.81E-6)

.MODEL RP+ RES (R=1.0 TC1=1.06E-3)

.MODEL DIOPIN1 D (IS=1E-25 RS=3.5E3 BV=6.2 IBV=1E-5)

.MODEL DIOPIN2 D (IS=2E-16 RS=450 CJO=892E-15 M=0.4 VJ=0.6)

.MODEL DIOCAP D (IS=1E-25 RS=310 BV=5.65 IBV=1E-5)

.MODEL DIOZEN D (IS=1E-25 RS=220 BV=5.95 IBV=1E-5)

.MODEL DRES200R D (CJO=5E-14, M=0.44, VJ=0.6, BV=18, IBV=1E-5, RS=150)

.MODEL DRES1K D (CJO=1E-13, M=0.44, VJ=0.6, BV=18, IBV=1E-5, RS=150)

.MODEL DRES5K D (CJO=2E-13, M=0.44, VJ=0.6, BV=18, IBV=1E-5, RS=150)

.MODEL DRES10K D (CJO=18E-14, M=0.44, VJ=0.6, BV=18, IBV=1E-5, RS=150)
**Power supplies
Vcc 18 0 DC +5
Vee 2 0 DC -5
*VinD+ 20 0 AC 10mV 0 
VinD+ 20 0 SIN 0 10mV 10k
VinD- 14 0 AC 0mV 0
*VinAB 13 0 AC 10mV 0

**jumpers
VaD- 17 19 DC 0
VaD+ 16 15 DC 0

**resistors
Rprobe 15 0 1Meg
R1 18 26 35.2k
*Rpa 18 19 15k
*Rpb 18 15 15k
*RA 8 9 32k  
*RB 9 10 18k
*R6 5 8 10k 
*R7 4 2 820

*** TOP LEVEL FACET: 2X1-LAYOUT{SCH}
QNODE267 15 14 22 2 SNPN_911
QNODE268 16 17 18 2 SPNP_911 0.5
QNODE257 16 17 18 2 SPNP_911 0.5
RNODE249 23 22 RP- 1K
RNODE232 28 25 RP- 1K
RNODE231 29 27 RP- 1K
RNODE229 2 29 RP- 1K
RNODE228 2 28 RP- 1K
QNODE219 23 26 25 2 SNPN_911
QNODE217 26 26 27 2 SNPN_911
*QNODE269 5 7 4 2 LNPN_911
*QNODE208 5 7 4 2 LNPN_911
*QNODE183 5 8 7 2 SNPN_911
*QNODE179 8 9 10 2 SNPN_911
*QNODE270 6 10 4 2 SPNP_911 0.5
*QNODE88 6 10 4 2 SPNP_911 0.5
*QNODE80 10 13 12 2 SNPN_911
*QNODE271 4 6 2 2 LNPN_911
*QNODE72 4 6 2 2 LNPN_911
RNODE24 23 21 RP- 1K
QNODE272 17 17 18 2 SPNP_911 0.5
QNODE16 17 17 18 2 SPNP_911 0.5
QNODE9 19 20 21 2 SNPN_911

*analysis request
*.AC DEC 100 1 1G
*.TRAN .1us 500us
.DC VinD+ -5 5 .1
.Probe
.END
